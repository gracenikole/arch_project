module fp_adder (srcA, srcB);
input [31:0] srcA;
input [31:0] srcB;

output [31:0] result;
output [3:0] ALUFlags;

wire N, Z, C, V;



endmodule //fp_adder