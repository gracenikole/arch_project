module fp_adder (
  
);

endmodule //fp_adder