// vim: set expandtab:

module condcheck (
    Cond,
    Flags,
    CondEx
);
    input wire [3:0] Cond;
    input wire [3:0] Flags;
    output wire CondEx;

    // ADD CODE HERE
endmodule
